parameter XY_SELECT_HL = 0;
parameter XY_SELECT_IX = 1;
parameter XY_SELECT_IY = 2;